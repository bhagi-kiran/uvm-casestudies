module add(add_if aif);

 assign aif.y = aif.a + aif.b;
endmodule
